`include "ahb_lite_slave.svp"
